module adjustment(
    
)